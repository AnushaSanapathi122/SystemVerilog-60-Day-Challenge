// Day 01: Introduction to SystemVerilog
// Simple hello program

module hello_systemverilog;
  initial begin
    $display("Hello SystemVerilog!");
    $display("Yahoooo!!!!.... Today(27-01-2025) I am Starting 60day system verilog challange");
  end
endmodule
